library verilog;
use verilog.vl_types.all;
entity risc_v32i_vlg_vec_tst is
end risc_v32i_vlg_vec_tst;
