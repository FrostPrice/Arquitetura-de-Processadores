library verilog;
use verilog.vl_types.all;
entity mux21_1b_vlg_vec_tst is
end mux21_1b_vlg_vec_tst;
