library verilog;
use verilog.vl_types.all;
entity add_sub_vlg_vec_tst is
end add_sub_vlg_vec_tst;
