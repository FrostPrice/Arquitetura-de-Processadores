library verilog;
use verilog.vl_types.all;
entity mux21_1b_vlg_check_tst is
    port(
        o_S             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux21_1b_vlg_check_tst;
